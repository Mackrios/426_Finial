library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity instruction_memory is
  port(
    address     : in  unsigned(15 downto 0);
    instruction : out unsigned(15 downto 0)
  );
end entity;

architecture rtl of instruction_memory is
  type mem_array is array(0 to 255) of unsigned(15 downto 0);


  
  
  
  signal mem : mem_array := (

    -- 0x00: addi r6, r6, -1
    -- [0011][110][110][111111]
    0  => x"3dbe",

    -- 0x02: addi r6, r6, -1
    -- [0011][110][110][111111]
    1  => x"3dbe",

    -- 0x04: addi r6, r6, -1
    -- [0011][110][110][111111]
    2  => x"3dbe",
    
    --3 => x"0000",
    
    --lw r1 r2 0 
    3 => x"1440",
    
    --addi r1 r1 -1
    4 => x"327f", 
    
    --5 => x"327f"


--    -- ============================================================
--    -- WHILE LOOP START (Address 0x00)
--    -- ============================================================

--    -- 0x00: addi r6, r6, -1
--    -- [0011][110][110][111111]
--    0  => x"04C8",

--    -- 0x02: lw r4, 0(r5)
--    -- [0001][101][100][000000]
--    1  => x"1B00",

--    -- 0x04: sub r7, r7, r7
--    -- [0000][111][111][111][001]
--    2  => x"0FF9",

--    -- 0x06: lw r7, 8(r7)
--    -- [0001][111][111][001000]
--    3  => x"1FE8",

--    -- 0x08: bgt r4, r7, +6
--    -- [0101][100][111][000110]
--    4  => x"59C6",

--    -- ============================================================
--    -- ELSE BRANCH (Address 0x0A)
--    -- ============================================================

--    -- 0x0A: sll r2, r2, 2
--    -- [0000][010][010][010][010]
--    5  => x"0492",

--    -- 0x0C: xor r3, r3, r2
--    -- [0000][011][010][011][111]
--    6  => x"069F",

--    -- 0x0E: lw r7, 10(r7)
--    -- [0001][111][111][001010]
--    7  => x"1FEA",

--    -- 0x10: sw r7, 0(r5)
--    -- [0010][101][111][000000]
--    8  => x"2BC0",

--    -- 0x12: j 0x20
--    -- [1000][000000100000]
--    9  => x"8020",

--    -- ============================================================
--    -- THEN BRANCH (Address 0x14)
--    -- ============================================================

--    -- 0x14: srl r0, r0, 3
--    -- [0000][000][000][000][011]   (shamt=3)
--    10 => x"0003",

--    -- 0x16: or r1, r1, r0
--    -- [0000][001][000][001][011]
--    11 => x"020B",

--    -- 0x18: sub r7, r7, r7
--    -- same encoding as before
--    12 => x"0FF9",

--    -- 0x1A: lw r7, 12(r7)
--    -- [0001][111][111][001100]
--    13 => x"1FEC",

--    -- 0x1C: sw r7, 0(r5)
--    -- [0010][101][111][000000]
--    14 => x"2BC0",

--    -- 0x1E: j 0x20
--    -- [1000][000000100000]
--    15 => x"8020",

--    -- ============================================================
--    -- ENDIF (Address 0x20)
--    -- ============================================================

--    -- 0x20: addi r5, r5, 2
--    -- [0011][101][101][000010]
--    16 => x"3B42",

--    -- 0x22: sub r7, r7, r7
--    17 => x"0FF9",

--    -- 0x24: bgt r6, r7, -18
--    -- imm(-18) = 101110
--    -- [0101][110][111][101110]
--    18 => x"5DEE",

--    -- ============================================================
--    -- RETURN / HALT (Address 0x26)
--    -- ============================================================

--    -- 0x26: j 0x26 (infinite loop)
--    -- [1000][000000100110]
--    19 => x"8026",

    others => (others => '0')
);

  
begin
  -- Word addressing: PC increments by 2 (byte addresses)
  instruction <= mem(to_integer(address(7 downto 1)));
end architecture;